
`timescale 1ns/1ps  
module SARSA_WInd_e8 (
input [1:0] A,
input [1:0] B,
output [3:0] P);

        // Generación de productos parciales
 wire pp0 = ((A[0]) & (B[0]));
 wire pp1 = ((1) & (B[1]));
 wire pp2 = ((A[1]) & (1));

    // Suma de productos parciales
wire [1:0] columna2 = pp1 + pp2;
wire [1:0] columna1 = pp0;


reg [3:0] corrected;
wire [3:0] rawP=(columna2 << 1) + (columna1 << 0); 

always @(*) begin
    case ({A,B})
      4'b1111: corrected = 4'd9; // ejemplo: A=0,B=3 => producto 0*3=0 (ajustar según necesidad)
      default: corrected = rawP;
    endcase
  end
assign P = corrected;
endmodule
