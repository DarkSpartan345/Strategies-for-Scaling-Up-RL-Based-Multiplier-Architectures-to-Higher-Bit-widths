
`timescale 1ns/1ps  
module SarsaNStepsRuido_e9 (
input [1:0] A,
input [1:0] B,
output [3:0] P);

        // Generación de productos parciales
 wire pp0 = ((A[1]) & (B[1]));
 wire pp1 = ((A[0]) & (1));
 wire pp2 = ((A[1]) & (B[0]));

    // Suma de productos parciales
wire [1:0] columna3 = pp0;
wire [1:0] columna2 = pp1 + pp2;
assign P = (columna3 << 2) + (columna2 << 1);
endmodule
